`timescale 1ns/100ps
module circ8(in0, in1, o0);
  input in0;
  input in1;

  output o0;
 
  and g5 (o0,in0,in1);
  
endmodule
